`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:56:40 03/03/2015 
// Design Name: 
// Module Name:    yx_cpu_mips16e 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module yx_cpu_mips16e(clk, rst);
	 
parameter word_size = 16;//the set_bits of cpu

input clk, rst;

//processing_unit
//M1_processing_unit ();
//control_unit
//M2_control_unit ();
//memory_unit
//M0_memory_unit ();

endmodule
